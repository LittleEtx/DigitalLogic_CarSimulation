`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/12/09 13:58:31
// Design Name: 
// Module Name: Engine
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Engine(
    input clk,
    input power_on,
    input power_off,
    input model_select,
    input throttle,
    input clutch,
    input brake,
    input reverse,
    input right,
    input left,
    input front_detector,
    input left_detector,
    input back_detector,
    input right_detector
    );
endmodule

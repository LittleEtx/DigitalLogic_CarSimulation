`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/12/09 14:10:53
// Design Name: 
// Module Name: semi_command
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module semi_command(
    input [1:0]state,
    input turn_left,
    input turn_right,
    input go_straight,
    output [1:0]cur,
    output clockwise
    );
endmodule

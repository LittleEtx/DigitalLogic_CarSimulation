`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/12/09 14:08:00
// Design Name: 
// Module Name: semi_state
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module semi_state(
    input [1:0]state,
    input front_detector,
    input back_detector,
    input left_detector,
    input right_detector,
    input clk,
    output [1:0]cur
    );



    
endmodule
